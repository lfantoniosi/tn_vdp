--
-- F18A
--   A pin-compatible enhanced replacement for the TMS9918A VDP family.
--   https://dnotq.io
--

-- Released under the 3-Clause BSD License:
--
-- Copyright 2011-2018 Matthew Hagerty (matthew <at> dnotq <dot> io)
--
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions are met:
--
-- 1. Redistributions of source code must retain the above copyright notice,
-- this list of conditions and the following disclaimer.
--
-- 2. Redistributions in binary form must reproduce the above copyright
-- notice, this list of conditions and the following disclaimer in the
-- documentation and/or other materials provided with the distribution.
--
-- 3. Neither the name of the copyright holder nor the names of its
-- contributors may be used to endorse or promote products derived from this
-- software without specific prior written permission.
--
-- THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
-- AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
-- IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE
-- ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE
-- LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR
-- CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF
-- SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS
-- INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN
-- CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE
-- POSSIBILITY OF SUCH DAMAGE.

-- Version history.  See README.md for details.
--
--   V1.9 Dec 31, 2018
--   V1.8 Aug 24, 2016
--   V1.7 Jan  1, 2016
--   V1.6 May  3, 2014 .. Apr 26, 2015
--   V1.5 Jul 23, 2013
--   V1.4 Mar 20, 2013 .. Apr 26, 2013
--   V1.3 Jul 26, 2012, Release firmware

-- The on-board 16K VRAM.  Initialized with font pattern and name table data
-- that will display the F18A power-on screen.  This allows the F18A to produce
-- a display even when there is no host CPU and helps troubleshooting.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity f18a_single_port_ram is
   port (
      clk   : in  std_logic;
      we    : in  std_logic;
      addr  : in  std_logic_vector(0 to 13);
      addr2 : in  std_logic_vector(0 to 13);
      din   : in  std_logic_vector(0 to 7);
      dout  : out std_logic_vector(0 to 7);
      dout2 : out std_logic_vector(0 to 7)
      );
end f18a_single_port_ram;

architecture rtl of f18a_single_port_ram is

   -- Initialize the VRAM with patterns for a font and credits / version information on the screen.
   type ram_t is array (0 to 16383) of std_logic_vector(0 to 7);
   signal ram : ram_t :=
   ( --  Comments on this line identify the version bytes --->                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       V     1     .     9                                                                             C     2     0     1     2     -     2     0     1     8
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"80",x"80",x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"81",x"81",x"00",x"00",x"03",x"03",x"03",x"03",x"00",x"00",x"00",x"00",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"00",x"00",x"C0",x"C0",x"E0",x"0F",x"0F",x"07",x"00",x"00",x"81",x"81",x"81",x"81",x"81",x"81",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"C0",x"C0",x"C0",x"E0",x"E0",x"00",x"00",x"00",x"00",x"80",x"80",x"80",x"C0",x"00",x"00",x"E0",x"C0",x"C0",x"C0",x"80",x"81",x"00",x"00",x"70",x"70",x"0F",x"0F",x"0F",x"0F",x"00",x"00",x"00",x"00",x"00",x"00",x"C1",x"C0",x"00",x"00",x"C0",x"0F",x"03",x"01",x"00",x"80",x"00",x"00",x"01",x"01",x"01",x"01",x"01",x"81",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"07",x"00",x"00",x"03",x"01",x"00",x"00",x"80",x"E0",x"00",x"00",x"00",x"00",x"80",x"80",x"C0",x"C0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"81",x"81",x"81",x"81",x"81",x"81",x"81",x"81",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"07",x"03",x"01",x"01",x"80",x"C0",x"C0",x"E0",x"81",x"81",x"81",x"81",x"81",x"81",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"E0",x"E0",x"E0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E0",x"0F",x"0F",x"0F",x"07",x"07",x"03",x"03",x"C0",x"C0",x"E0",x"E0",x"1E",x"0E",x"0E",x"0C",x"81",x"01",x"03",x"03",x"03",x"07",x"07",x"07",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"81",x"81",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"07",x"07",x"07",x"07",x"07",x"07",x"00",x"00",x"0F",x"0F",x"0F",x"E0",x"E0",x"80",x"00",x"00",x"C0",x"C0",x"C0",x"C0",x"C0",x"80",x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"81",x"81",x"81",x"81",x"81",x"81",x"81",x"81",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"E0",x"0F",x"07",x"07",x"03",x"03",x"01",x"00",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"E0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"01",x"01",x"01",x"00",x"00",x"00",x"00",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"80",x"0F",x"0F",x"E0",x"E0",x"E0",x"C0",x"C0",x"C0",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"C0",x"C0",x"C0",x"C0",x"C0",x"C1",x"00",x"00",x"E0",x"E0",x"E0",x"C0",x"80",x"00",x"01",x"03",x"C1",x"C1",x"81",x"81",x"01",x"01",x"01",x"01",x"00",x"00",x"07",x"07",x"07",x"07",x"07",x"07",x"01",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"80",x"80",x"80",x"81",x"81",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"C0",x"C0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"81",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"0F",x"0F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0F",x"C0",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E0",x"E0",x"E0",x"E0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3C",x"42",x"5A",x"81",x"5A",x"66",x"42",x"3C",x"3C",x"81",x"24",x"00",x"00",x"24",x"66",x"3C",x"6C",x"01",x"01",x"01",x"83",x"38",x"10",x"00",x"10",x"38",x"83",x"01",x"83",x"38",x"10",x"00",x"10",x"38",x"54",x"01",x"54",x"10",x"38",x"00",x"10",x"38",x"83",x"01",x"01",x"10",x"38",x"00",x"00",x"00",x"00",x"30",x"30",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"00",x"00",x"00",x"38",x"44",x"82",x"82",x"82",x"44",x"38",x"00",x"38",x"44",x"82",x"82",x"82",x"44",x"38",x"00",x"0F",x"03",x"05",x"86",x"88",x"88",x"88",x"70",x"38",x"44",x"44",x"44",x"38",x"10",x"83",x"10",x"30",x"28",x"24",x"24",x"28",x"20",x"E0",x"C0",x"3C",x"24",x"3C",x"24",x"24",x"1B",x"23",x"18",x"10",x"54",x"38",x"11",x"38",x"54",x"10",x"00",x"10",x"10",x"10",x"83",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"0F",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"E0",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E0",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"0F",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"E0",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"0F",x"00",x"00",x"00",x"00",x"81",x"42",x"24",x"18",x"18",x"24",x"42",x"81",x"01",x"02",x"04",x"08",x"10",x"20",x"40",x"80",x"80",x"40",x"20",x"10",x"08",x"04",x"02",x"01",x"00",x"10",x"10",x"00",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"00",x"00",x"20",x"00",x"50",x"50",x"50",x"00",x"00",x"00",x"00",x"00",x"50",x"50",x"07",x"50",x"07",x"50",x"50",x"00",x"20",x"78",x"A0",x"70",x"28",x"0F",x"20",x"00",x"C0",x"C8",x"10",x"20",x"40",x"98",x"18",x"00",x"40",x"A0",x"40",x"A8",x"90",x"98",x"60",x"00",x"10",x"20",x"40",x"00",x"00",x"00",x"00",x"00",x"10",x"20",x"40",x"40",x"40",x"20",x"10",x"00",x"40",x"20",x"10",x"10",x"10",x"20",x"40",x"00",x"20",x"A8",x"70",x"20",x"70",x"A8",x"20",x"00",x"00",x"20",x"20",x"07",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"40",x"00",x"00",x"00",x"78",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"60",x"60",x"00",x"00",x"00",x"08",x"10",x"20",x"40",x"80",x"00",x"70",x"88",x"98",x"A8",x"C8",x"88",x"70",x"00",x"20",x"60",x"A0",x"20",x"20",x"20",x"07",x"00",x"70",x"88",x"08",x"10",x"60",x"80",x"07",x"00",x"70",x"88",x"08",x"30",x"08",x"88",x"70",x"00",x"10",x"30",x"50",x"90",x"07",x"10",x"10",x"00",x"07",x"80",x"E0",x"10",x"08",x"10",x"E0",x"00",x"30",x"40",x"80",x"0F",x"88",x"88",x"70",x"00",x"07",x"88",x"10",x"20",x"20",x"20",x"20",x"00",x"70",x"88",x"88",x"70",x"88",x"88",x"70",x"00",x"70",x"88",x"88",x"78",x"08",x"10",x"60",x"00",x"00",x"00",x"20",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"20",x"20",x"40",x"18",x"30",x"60",x"C0",x"60",x"30",x"18",x"00",x"00",x"00",x"07",x"00",x"07",x"00",x"00",x"00",x"C0",x"60",x"30",x"18",x"30",x"60",x"C0",x"00",x"70",x"88",x"08",x"10",x"20",x"00",x"20",x"00",x"70",x"88",x"08",x"68",x"A8",x"A8",x"70",x"00",x"20",x"50",x"88",x"88",x"07",x"88",x"88",x"00",x"0F",x"48",x"48",x"70",x"48",x"48",x"0F",x"00",x"30",x"48",x"80",x"80",x"80",x"48",x"30",x"00",x"E0",x"50",x"48",x"48",x"48",x"50",x"E0",x"00",x"07",x"80",x"80",x"0F",x"80",x"80",x"07",x"00",x"07",x"80",x"80",x"0F",x"80",x"80",x"80",x"00",x"70",x"88",x"80",x"47",x"88",x"88",x"70",x"00",x"88",x"88",x"88",x"07",x"88",x"88",x"88",x"00",x"70",x"20",x"20",x"20",x"20",x"20",x"70",x"00",x"38",x"10",x"10",x"10",x"90",x"90",x"60",x"00",x"88",x"90",x"A0",x"C0",x"A0",x"90",x"88",x"00",x"80",x"80",x"80",x"80",x"80",x"80",x"07",x"00",x"88",x"27",x"A8",x"A8",x"88",x"88",x"88",x"00",x"88",x"C8",x"C8",x"A8",x"98",x"98",x"88",x"00",x"70",x"88",x"88",x"88",x"88",x"88",x"70",x"00",x"0F",x"88",x"88",x"0F",x"80",x"80",x"80",x"00",x"70",x"88",x"88",x"88",x"A8",x"90",x"68",x"00",x"0F",x"88",x"88",x"0F",x"A0",x"90",x"88",x"00",x"70",x"88",x"80",x"70",x"08",x"88",x"70",x"00",x"07",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"88",x"88",x"88",x"88",x"88",x"88",x"70",x"00",x"88",x"88",x"88",x"88",x"50",x"50",x"20",x"00",x"88",x"88",x"88",x"A8",x"A8",x"27",x"88",x"00",x"88",x"88",x"50",x"20",x"50",x"88",x"88",x"00",x"88",x"88",x"88",x"70",x"20",x"20",x"20",x"00",x"07",x"08",x"10",x"20",x"40",x"80",x"07",x"00",x"70",x"40",x"40",x"40",x"40",x"40",x"70",x"00",x"00",x"00",x"80",x"40",x"20",x"10",x"08",x"00",x"70",x"10",x"10",x"10",x"10",x"10",x"70",x"00",x"20",x"50",x"88",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"00",x"40",x"20",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"70",x"08",x"78",x"88",x"78",x"00",x"80",x"80",x"B0",x"C8",x"88",x"C8",x"B0",x"00",x"00",x"00",x"70",x"88",x"80",x"88",x"70",x"00",x"08",x"08",x"68",x"98",x"88",x"98",x"68",x"00",x"00",x"00",x"70",x"88",x"07",x"80",x"70",x"00",x"10",x"28",x"20",x"07",x"20",x"20",x"20",x"00",x"00",x"00",x"68",x"98",x"98",x"68",x"08",x"70",x"80",x"80",x"0F",x"88",x"88",x"88",x"88",x"00",x"20",x"00",x"60",x"20",x"20",x"20",x"70",x"00",x"10",x"00",x"30",x"10",x"10",x"10",x"90",x"60",x"40",x"40",x"48",x"50",x"60",x"50",x"48",x"00",x"60",x"20",x"20",x"20",x"20",x"20",x"70",x"00",x"00",x"00",x"D0",x"A8",x"A8",x"A8",x"A8",x"00",x"00",x"00",x"B0",x"C8",x"88",x"88",x"88",x"00",x"00",x"00",x"70",x"88",x"88",x"88",x"70",x"00",x"00",x"00",x"B0",x"C8",x"C8",x"B0",x"80",x"80",x"00",x"00",x"68",x"98",x"98",x"68",x"08",x"08",x"00",x"00",x"B0",x"C8",x"80",x"80",x"80",x"00",x"00",x"00",x"78",x"80",x"0F",x"08",x"0F",x"00",x"40",x"40",x"0F",x"40",x"40",x"48",x"30",x"00",x"00",x"00",x"90",x"90",x"90",x"90",x"68",x"00",x"00",x"00",x"88",x"88",x"88",x"50",x"20",x"00",x"00",x"00",x"88",x"A8",x"A8",x"A8",x"50",x"00",x"00",x"00",x"88",x"50",x"20",x"50",x"88",x"00",x"00",x"00",x"88",x"88",x"98",x"68",x"08",x"70",x"00",x"00",x"07",x"10",x"20",x"40",x"07",x"00",x"18",x"20",x"20",x"40",x"20",x"20",x"18",x"00",x"20",x"20",x"20",x"00",x"20",x"20",x"20",x"00",x"C0",x"20",x"20",x"10",x"20",x"20",x"C0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"70",x"88",x"80",x"80",x"88",x"70",x"20",x"60",x"90",x"00",x"00",x"90",x"90",x"90",x"68",x"00",x"10",x"20",x"70",x"88",x"07",x"80",x"70",x"00",x"20",x"50",x"70",x"08",x"78",x"88",x"78",x"00",x"48",x"00",x"70",x"08",x"78",x"88",x"78",x"00",x"20",x"10",x"70",x"08",x"78",x"88",x"78",x"00",x"20",x"00",x"70",x"08",x"78",x"88",x"78",x"00",x"00",x"70",x"80",x"80",x"80",x"70",x"10",x"60",x"20",x"50",x"70",x"88",x"07",x"80",x"70",x"00",x"50",x"00",x"70",x"88",x"07",x"80",x"70",x"00",x"20",x"10",x"70",x"88",x"07",x"80",x"70",x"00",x"50",x"00",x"00",x"60",x"20",x"20",x"70",x"00",x"20",x"50",x"00",x"60",x"20",x"20",x"70",x"00",x"40",x"20",x"00",x"60",x"20",x"20",x"70",x"00",x"50",x"00",x"20",x"50",x"88",x"07",x"88",x"00",x"20",x"00",x"20",x"50",x"88",x"07",x"88",x"00",x"10",x"20",x"07",x"80",x"0F",x"80",x"07",x"00",x"00",x"00",x"6C",x"12",x"81",x"90",x"91",x"00",x"C1",x"50",x"90",x"63",x"0F",x"90",x"61",x"00",x"60",x"90",x"00",x"60",x"90",x"90",x"60",x"00",x"90",x"00",x"00",x"60",x"90",x"90",x"60",x"00",x"40",x"20",x"00",x"60",x"90",x"90",x"60",x"00",x"40",x"A0",x"00",x"A0",x"A0",x"A0",x"50",x"00",x"40",x"20",x"00",x"A0",x"A0",x"A0",x"50",x"00",x"90",x"00",x"90",x"90",x"B0",x"50",x"10",x"E0",x"50",x"00",x"70",x"88",x"88",x"88",x"70",x"00",x"50",x"00",x"88",x"88",x"88",x"88",x"70",x"00",x"20",x"20",x"78",x"80",x"80",x"78",x"20",x"20",x"18",x"24",x"20",x"07",x"20",x"1D",x"5C",x"00",x"88",x"50",x"20",x"07",x"20",x"07",x"20",x"00",x"C0",x"A0",x"A0",x"C8",x"63",x"88",x"88",x"8C",x"18",x"20",x"20",x"07",x"20",x"20",x"20",x"40",x"10",x"20",x"70",x"08",x"78",x"88",x"78",x"00",x"10",x"20",x"00",x"60",x"20",x"20",x"70",x"00",x"20",x"40",x"00",x"60",x"90",x"90",x"60",x"00",x"20",x"40",x"00",x"90",x"90",x"90",x"68",x"00",x"50",x"A0",x"00",x"A0",x"D0",x"90",x"90",x"00",x"28",x"50",x"00",x"C8",x"A8",x"98",x"88",x"00",x"00",x"70",x"08",x"78",x"88",x"78",x"00",x"07",x"00",x"60",x"90",x"90",x"90",x"60",x"00",x"0F",x"20",x"00",x"20",x"40",x"80",x"88",x"70",x"00",x"00",x"00",x"00",x"07",x"80",x"80",x"00",x"00",x"00",x"00",x"00",x"07",x"08",x"08",x"00",x"00",x"84",x"88",x"90",x"A8",x"54",x"84",x"08",x"1C",x"84",x"88",x"90",x"A8",x"58",x"A8",x"3C",x"08",x"20",x"00",x"00",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"24",x"48",x"90",x"48",x"24",x"00",x"00",x"00",x"90",x"48",x"24",x"48",x"90",x"00",x"28",x"50",x"20",x"50",x"88",x"07",x"88",x"00",x"28",x"50",x"70",x"08",x"78",x"88",x"78",x"00",x"28",x"50",x"00",x"70",x"20",x"20",x"70",x"00",x"28",x"50",x"00",x"20",x"20",x"20",x"70",x"00",x"28",x"50",x"00",x"70",x"88",x"88",x"70",x"00",x"50",x"A0",x"00",x"60",x"90",x"90",x"60",x"00",x"28",x"50",x"00",x"88",x"88",x"88",x"70",x"00",x"50",x"A0",x"00",x"A0",x"A0",x"A0",x"50",x"00",x"03",x"48",x"48",x"48",x"17",x"08",x"50",x"20",x"00",x"50",x"00",x"50",x"50",x"50",x"10",x"20",x"C0",x"44",x"C8",x"54",x"13",x"54",x"61",x"04",x"10",x"A8",x"40",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"50",x"88",x"50",x"20",x"00",x"00",x"88",x"10",x"20",x"40",x"80",x"28",x"00",x"00",x"83",x"A8",x"A8",x"68",x"28",x"28",x"28",x"00",x"38",x"40",x"30",x"48",x"48",x"30",x"08",x"70",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3C",x"3C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"11",x"22",x"44",x"88",x"11",x"22",x"44",x"88",x"88",x"44",x"22",x"11",x"88",x"44",x"22",x"11",x"01",x"83",x"38",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"38",x"83",x"01",x"80",x"C0",x"E0",x"0F",x"E0",x"C0",x"80",x"00",x"01",x"03",x"07",x"0F",x"07",x"03",x"01",x"00",x"00",x"81",x"3C",x"18",x"18",x"3C",x"81",x"00",x"81",x"3C",x"18",x"00",x"00",x"18",x"3C",x"81",x"0F",x"0F",x"0F",x"0F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0F",x"0F",x"0F",x"0F",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"00",x"20",x"20",x"50",x"50",x"88",x"07",x"00",x"20",x"20",x"70",x"20",x"70",x"20",x"20",x"00",x"00",x"00",x"00",x"50",x"88",x"A8",x"50",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3C",x"42",x"5A",x"81",x"5A",x"66",x"42",x"3C",x"3C",x"81",x"24",x"00",x"00",x"24",x"66",x"3C",x"6C",x"01",x"01",x"01",x"83",x"38",x"10",x"00",x"10",x"38",x"83",x"01",x"83",x"38",x"10",x"00",x"10",x"38",x"54",x"01",x"54",x"10",x"38",x"00",x"10",x"38",x"83",x"01",x"01",x"10",x"38",x"00",x"00",x"00",x"00",x"30",x"30",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"00",x"00",x"00",x"38",x"44",x"82",x"82",x"82",x"44",x"38",x"00",x"38",x"44",x"82",x"82",x"82",x"44",x"38",x"00",x"0F",x"03",x"05",x"86",x"88",x"88",x"88",x"70",x"38",x"44",x"44",x"44",x"38",x"10",x"83",x"10",x"30",x"28",x"24",x"24",x"28",x"20",x"E0",x"C0",x"3C",x"24",x"3C",x"24",x"24",x"1B",x"23",x"18",x"10",x"54",x"38",x"11",x"38",x"54",x"10",x"00",x"10",x"10",x"10",x"83",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"0F",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"E0",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E0",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"0F",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"E0",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"0F",x"00",x"00",x"00",x"00",x"81",x"42",x"24",x"18",x"18",x"24",x"42",x"81",x"01",x"02",x"04",x"08",x"10",x"20",x"40",x"80",x"80",x"40",x"20",x"10",x"08",x"04",x"02",x"01",x"00",x"10",x"10",x"00",x"10",x"10",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"01",x"02",x"03",x"04",x"05",x"06",x"07",x"08",x"09",x"0A",x"0B",x"0C",x"0D",x"0E",x"0F",x"10",x"11",x"12",x"13",x"14",x"15",x"16",x"17",x"18",x"19",x"1A",x"1B",x"1C",x"1D",x"1E",x"1F",x"20",x"21",x"22",x"23",x"24",x"25",x"26",x"27",x"28",x"29",x"2A",x"2B",x"2C",x"2D",x"2E",x"2F",x"30",x"31",x"32",x"33",x"34",x"35",x"36",x"37",x"38",x"39",x"3A",x"3B",x"3C",x"3D",x"3E",x"3F",x"40",x"41",x"42",x"43",x"44",x"45",x"46",x"47",x"48",x"49",x"4A",x"4B",x"4C",x"4D",x"4E",x"4F",x"50",x"51",x"52",x"53",x"54",x"55",x"56",x"57",x"58",x"59",x"5A",x"5B",x"5C",x"5D",x"5E",x"5F",x"60",x"61",x"62",x"63",x"64",x"65",x"66",x"67",x"68",x"69",x"6A",x"6B",x"6C",x"6D",x"6E",x"6F",x"70",x"71",x"72",x"73",x"74",x"75",x"76",x"77",x"78",x"79",x"7A",x"7B",x"7C",x"7D",x"7E",x"7F",x"80",x"81",x"82",x"83",x"84",x"85",x"86",x"87",x"88",x"89",x"8A",x"8B",x"8C",x"8D",x"8E",x"8F",x"90",x"91",x"92",x"93",x"94",x"95",x"96",x"97",x"98",x"99",x"9A",x"9B",x"9C",x"9D",x"9E",x"9F",x"A0",x"A1",x"A2",x"A3",x"A4",x"A5",x"A6",x"A7",x"A8",x"A9",x"AA",x"AB",x"AC",x"AD",x"AE",x"AF",x"B0",x"B1",x"B2",x"B3",x"B4",x"B5",x"B6",x"B7",x"B8",x"B9",x"BA",x"BB",x"BC",x"BD",x"BE",x"BF",x"C0",x"C1",x"C2",x"C3",x"C4",x"C5",x"C6",x"C7",x"C8",x"C9",x"CA",x"CB",x"CC",x"CD",x"CE",x"CF",x"D0",x"D1",x"D2",x"D3",x"D4",x"D5",x"D6",x"D7",x"D8",x"D9",x"DA",x"DB",x"DC",x"DD",x"DE",x"DF",x"E0",x"E1",x"E2",x"E3",x"E4",x"E5",x"E6",x"E7",x"E8",x"E9",x"EA",x"EB",x"EC",x"ED",x"EE",x"EF",x"F0",x"F1",x"F2",x"F3",x"F4",x"F5",x"F6",x"F7",x"F8",x"F9",x"FA",x"FB",x"FC",x"FD",x"FE",x"FF",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"2D",x"2D",x"2D",x"2D",x"2D",x"2D",x"2D",x"2D",x"2D",x"2D",x"2D",x"2D",x"2D",x"2D",x"2D",x"2D",x"2D",x"2D",x"2D",x"2D",x"2D",x"2D",x"2D",x"2D",x"2D",x"2D",x"20",x"20",x"20",x"20",x"20",x"20",x"54",x"41",x"4E",x"47",x"20",x"4E",x"41",x"4E",x"4F",x"20",x"39",x"4B",x"20",x"20",x"54",x"4D",x"53",x"39",x"39",x"31",x"38",x"41",x"20",x"56",x"44",x"50",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"31",x"36",x"4B",x"42",x"20",x"56",x"52",x"41",x"4D",x"20",x"2D",x"20",x"48",x"44",x"4D",x"49",x"2F",x"41",x"55",x"44",x"49",x"4F",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"56",x"45",x"52",x"53",x"49",x"4F",x"4E",x"20",x"32",x"2E",x"30",x"30",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"2D",x"2D",x"2D",x"2D",x"2D",x"2D",x"2D",x"2D",x"2D",x"2D",x"2D",x"2D",x"2D",x"2D",x"2D",x"2D",x"2D",x"2D",x"2D",x"2D",x"2D",x"2D",x"2D",x"2D",x"2D",x"2D",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"01",x"02",x"03",x"04",x"05",x"06",x"07",x"08",x"09",x"0A",x"0B",x"0C",x"0D",x"0E",x"0F",x"10",x"11",x"12",x"13",x"14",x"15",x"16",x"17",x"18",x"19",x"1A",x"1B",x"1C",x"1D",x"1E",x"1F",x"20",x"21",x"22",x"23",x"24",x"25",x"26",x"27",x"28",x"29",x"2A",x"2B",x"2C",x"2D",x"2E",x"2F",x"30",x"31",x"32",x"33",x"34",x"35",x"36",x"37",x"38",x"39",x"3A",x"3B",x"3C",x"3D",x"3E",x"3F",x"40",x"41",x"42",x"43",x"44",x"45",x"46",x"47",x"48",x"49",x"4A",x"4B",x"4C",x"4D",x"4E",x"4F",x"50",x"51",x"52",x"53",x"54",x"55",x"56",x"57",x"58",x"59",x"5A",x"5B",x"5C",x"5D",x"5E",x"5F",x"60",x"61",x"62",x"63",x"64",x"65",x"66",x"67",x"68",x"69",x"6A",x"6B",x"6C",x"6D",x"6E",x"6F",x"70",x"71",x"72",x"73",x"74",x"75",x"76",x"77",x"78",x"79",x"7A",x"7B",x"7C",x"7D",x"7E",x"7F",x"80",x"81",x"82",x"83",x"84",x"85",x"86",x"87",x"88",x"89",x"8A",x"8B",x"8C",x"8D",x"8E",x"8F",x"90",x"91",x"92",x"93",x"94",x"95",x"96",x"97",x"98",x"99",x"9A",x"9B",x"9C",x"9D",x"9E",x"9F",x"A0",x"A1",x"A2",x"A3",x"A4",x"A5",x"A6",x"A7",x"A8",x"A9",x"AA",x"AB",x"AC",x"AD",x"AE",x"AF",x"B0",x"B1",x"B2",x"B3",x"B4",x"B5",x"B6",x"B7",x"B8",x"B9",x"BA",x"BB",x"BC",x"BD",x"BE",x"BF",x"C0",x"C1",x"C2",x"C3",x"C4",x"C5",x"C6",x"C7",x"C8",x"C9",x"CA",x"CB",x"CC",x"CD",x"CE",x"CF",x"D0",x"D1",x"D2",x"D3",x"D4",x"D5",x"D6",x"D7",x"D8",x"D9",x"DA",x"DB",x"DC",x"DD",x"DE",x"DF",x"E0",x"E1",x"E2",x"E3",x"E4",x"E5",x"E6",x"E7",x"E8",x"E9",x"EA",x"EB",x"EC",x"ED",x"EE",x"EF",x"F0",x"F1",x"F2",x"F3",x"F4",x"F5",x"F6",x"F7",x"F8",x"F9",x"FA",x"FB",x"FC",x"FD",x"FE",x"FF",x"D1",x"00",x"00",x"0F",x"D1",x"00",x"01",x"0F",x"D1",x"00",x"02",x"0F",x"D1",x"00",x"03",x"0F",x"D1",x"00",x"04",x"0F",x"D1",x"00",x"05",x"0F",x"D1",x"00",x"06",x"0F",x"D1",x"00",x"07",x"0F",x"D1",x"00",x"08",x"0F",x"D1",x"00",x"09",x"0F",x"D1",x"00",x"0A",x"0F",x"D1",x"00",x"0B",x"0F",x"D1",x"00",x"0C",x"0F",x"D1",x"00",x"0D",x"0F",x"D1",x"00",x"0E",x"0F",x"D1",x"00",x"0F",x"0F",x"D1",x"00",x"10",x"0F",x"D1",x"00",x"11",x"0F",x"D1",x"00",x"12",x"0F",x"D1",x"00",x"13",x"0F",x"D1",x"00",x"14",x"0F",x"D1",x"00",x"15",x"0F",x"D1",x"00",x"16",x"0F",x"D1",x"00",x"17",x"0F",x"D1",x"00",x"18",x"0F",x"D1",x"00",x"19",x"0F",x"D1",x"00",x"1A",x"0F",x"D1",x"00",x"1B",x"0F",x"D1",x"00",x"1C",x"0F",x"D1",x"00",x"1D",x"0F",x"D1",x"00",x"1E",x"0F",x"D1",x"00",x"1F",x"0F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0F",x"0F",x"0F",x"0F",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"0F",x"0F",x"00",x"00",x"0F",x"0F",x"0F",x"0F",x"00",x"00",x"00",x"00",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"00",x"00",x"F0",x"F0",x"F0",x"0F",x"0F",x"0F",x"00",x"00",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"00",x"00",x"00",x"00",x"F0",x"F0",x"F0",x"F0",x"00",x"00",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"00",x"00",x"0F",x"0F",x"F0",x"F0",x"F0",x"F0",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"F0",x"F0",x"00",x"00",x"F0",x"0F",x"0F",x"0F",x"FF",x"0F",x"00",x"00",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"0F",x"0F",x"00",x"00",x"0F",x"0F",x"FF",x"FF",x"0F",x"0F",x"00",x"00",x"00",x"00",x"F0",x"F0",x"F0",x"F0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"00",x"00",x"00",x"00",x"00",x"0F",x"0F",x"0F",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"0F",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"FF",x"FF",x"F0",x"F0",x"F0",x"0F",x"0F",x"0F",x"FF",x"FF",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",
x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"00",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"F0",x"F0",x"F0",x"F0",x"00",x"00",x"00",x"00",x"0F",x"0F",x"FF",x"FF",x"FF",x"FF",x"FF",x"0F",x"0F",x"0F",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"FF",x"FF",x"0F",x"0F",x"0F",x"0F",x"0F",x"FF",x"0F",x"0F",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"FF",x"FF",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"0F",x"0F",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"0F",x"0F",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"0F",x"0F",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"F0",x"F0",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"F0",x"F0",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"0F",x"F0",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"F0",x"F0",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"0F",x"0F",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"F0",x"F0",x"F0",x"F0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",
x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"F4",x"F4",x"4F",x"F4",x"4F",x"4F",x"F4",x"F4",x"F4",x"4F",x"4F",x"FF",x"FF",x"4F",x"F4",x"F4",x"F4",x"4F",x"4F",x"4F",x"4F",x"F4",x"F4",x"44",x"F4",x"F4",x"4F",x"4F",x"4F",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"4F",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"4F",x"4F",x"4F",x"F4",x"F4",x"44",x"44",x"44",x"44",x"F4",x"F4",x"44",x"44",x"44",x"FF",x"FF",x"FF",x"4F",x"4F",x"FF",x"FF",x"FF",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"FF",x"F4",x"F4",x"F4",x"4F",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"4F",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"4F",x"4F",x"F4",x"F4",x"F4",x"F4",x"4F",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"4F",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"FF",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"FF",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"4F",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"4F",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"FF",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"44",x"44",x"FF",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"4F",x"F4",x"F4",x"F4",x"F4",x"44",x"44",x"44",x"4F",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"4F",x"44",x"44",x"44",x"44",x"F4",x"F4",x"F4",x"4F",x"44",x"44",x"44",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"FF",x"F4",x"F4",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"F4",x"F4",x"F4",x"F4",x"44",x"44",x"F4",x"44",x"F4",x"F4",x"F4",x"44",x"44",x"44",x"44",x"44",x"F4",x"F4",x"4F",x"F4",x"4F",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"4F",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"44",x"44",x"44",x"44",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"44",x"F4",x"F4",x"4F",x"F4",x"F4",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"F4",x"F4",x"F4",x"44",x"44",x"44",x"F4",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"F4",x"F4",x"44",x"44",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"4F",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"4F",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"4F",x"F4",x"F4",x"44",x"4F",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"4F",x"F4",x"F4",x"F4",x"44",x"4F",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"44",x"44",x"F4",x"44",x"44",x"F4",x"44",x"44",x"44",x"44",x"F4",x"44",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"44",x"44",x"4F",x"44",x"4F",x"44",x"44",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"4F",x"F4",x"F4",x"44",x"4F",x"F4",x"F4",x"F4",x"F4",x"F4",x"4F",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"4F",x"F4",x"F4",x"4F",x"F4",x"F4",x"4F",x"44",x"4F",x"F4",x"F4",x"4F",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"4F",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"4F",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"4F",x"44",x"F4",x"4F",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"4F",x"F4",x"F4",x"4F",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"4F",x"F4",x"F4",x"4F",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"4F",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"4F",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"4F",x"F4",x"F4",x"F4",x"F4",x"F4",x"4F",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"44",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"4F",x"44",x"F4",x"F4",x"F4",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"44",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"44",x"44",x"F4",x"F4",x"4F",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"4F",x"F4",x"F4",x"F4",x"44",x"44",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"4F",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"44",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"44",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"44",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"44",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"44",x"44",x"F4",x"F4",x"4F",x"F4",x"4F",x"44",x"F4",x"F4",x"4F",x"F4",x"F4",x"F4",x"F4",x"44",x"44",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"44",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"44",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"44",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"44",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"44",x"4F",x"F4",x"F4",x"F4",x"4F",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"44",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"4F",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"4F",x"F4",x"F4",x"44",x"F4",x"44",x"F4",x"F4",x"4F",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"4F",x"F4",x"F4",x"44",x"F4",x"44",x"44",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"44",x"F4",x"F4",x"F4",x"4F",x"F4",x"44",x"F4",x"44",x"F4",x"F4",x"F4",x"4F",x"F4",x"44",x"F4",x"F4",x"4F",x"F4",x"4F",x"F4",x"4F",x"44",x"44",x"44",x"F4",x"F4",x"4F",x"F4",x"4F",x"44",x"4F",x"F4",x"F4",x"4F",x"4F",x"F4",x"4F",x"44",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"44",x"44",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"4F",x"F4",x"4F",x"F4",x"44",x"F4",x"F4",x"F4",x"4F",x"F4",x"4F",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"4F",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"4F",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"44",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"4F",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"4F",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"44",x"44",x"44",x"4F",x"F4",x"F4",x"44",x"44",x"44",x"44",x"44",x"4F",x"F4",x"F4",x"44",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"44",x"F4",x"F4",x"F4",x"F4",x"44",x"44",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"44",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"4F",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"44",x"4F",x"F4",x"F4",x"F4",x"4F",x"F4",x"F4",x"F4",x"44",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"4F",x"F4",x"4F",x"F4",x"F4",x"F4",x"F4",x"44",x"44",x"44",x"44",x"44",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"44",x"4F",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"44",x"44",x"44",x"44",x"44",x"FF",x"FF",x"4F",x"4F",x"4F",x"4F",x"F4",x"F4",x"F4",x"F4",x"44",x"44",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"F4",x"F4",x"44",x"44",x"44",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"44",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"4F",x"4F",x"F4",x"F4",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"F4",x"F4",x"4F",x"4F",x"F4",x"F4",x"F4",x"4F",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"FF",x"4F",x"F4",x"F4",x"F4",x"F4",x"4F",x"FF",x"F4",x"4F",x"4F",x"FF",x"FF",x"4F",x"4F",x"F4",x"4F",x"4F",x"4F",x"4F",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"4F",x"4F",x"4F",x"4F",x"F4",x"F4",x"4F",x"4F",x"F4",x"F4",x"4F",x"4F",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"4F",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"44",x"44",x"44",x"F4",x"F4",x"F4",x"F4",x"44",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"44",x"44",x"44",x"44",x"FF",x"FF",x"FF",x"FF",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"FF",x"FF",x"FF",x"FF",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"F4",x"F4",x"4F",x"F4",x"4F",x"4F",x"F4",x"F4",x"F4",x"4F",x"4F",x"FF",x"FF",x"4F",x"F4",x"F4",x"F4",x"4F",x"4F",x"4F",x"4F",x"F4",x"F4",x"44",x"F4",x"F4",x"4F",x"4F",x"4F",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"4F",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"4F",x"4F",x"4F",x"F4",x"F4",x"44",x"44",x"44",x"44",x"F4",x"F4",x"44",x"44",x"44",x"FF",x"FF",x"FF",x"4F",x"4F",x"FF",x"FF",x"FF",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"FF",x"F4",x"F4",x"F4",x"4F",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"4F",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"4F",x"4F",x"F4",x"F4",x"F4",x"F4",x"4F",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"F4",x"4F",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"FF",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"FF",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"4F",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"4F",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"FF",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"44",x"44",x"FF",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"4F",x"F4",x"F4",x"F4",x"F4",x"44",x"44",x"44",x"4F",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"4F",x"44",x"44",x"44",x"44",x"F4",x"F4",x"F4",x"4F",x"44",x"44",x"44",x"44",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"44",x"F4",x"F4",x"FF",x"F4",x"F4",x"44",x"44",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
);

begin
   -- Inferred read_first ram.
   process (clk)
   begin
      if rising_edge(clk) then
         dout <= ram(to_integer(unsigned(addr)));
         dout2 <= ram(to_integer(unsigned(addr2)));
         if we = '1' then
            ram(to_integer(unsigned(addr))) <= din;
         end if;
      end if;
   end process;

end rtl;
